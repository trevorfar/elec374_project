`timescale 1ns / 1ps

module booth_mul_32_tb;

reg signed [31:0] a;
reg signed [31:0] b;
wire signed [63:0] cout;

booth_mul_32 uut(.M_input(a), .Q_input(b), .Z(cout));
initial begin
		  a = 32'b0000_0000_0000_0000_0000_0000_0000_0100; b = 32'b0000_0000_0000_0000_0000_0000_0000_0011; 
		  #50;
		  a = 32'b0000_0000_0000_0000_0000_0000_0000_0100; b = 32'b1111_1111_1111_1111_1111_1111_1111_1101;
		  #50
		  a = 32'b1111_1111_1111_1111_1111_1111_1111_1100; b = 32'b1111_1111_1111_1111_1111_1111_1111_1101;
		  #50
		  a = 32'b0; b = 32'b1111_1111_1111_1111_1111_1111_1111_1101;
		  #50
		 $stop;
end
endmodule


