`timescale 1ns / 1ps


module or_32_bit_tb;
reg [31:0] a;
reg [31:0] b;
wire [31:0] z;

or_32_bit uut(.a(a), .b(b), .z(z));
initial begin
		  a = 32'b0000_0000_0000_0000_0000_0000_0000_0000; b = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
		  #50;
		  a = 32'b1111_1111_1111_1111_1111_1111_1111_1111; b = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
		  #50
		  a = 32'b1111_1111_1111_1111_1111_1111_1111_1100; b = 32'b1111_1111_1111_1111_1111_1111_1111_1101;
		  #50
		  a = 32'b1111; b = 32'b1111;
		  #50
		  a = 32'b0001; b = 32'b0001;
		  #50
		  a = 32'b0101; b = 32'b1010;
		 $stop;
end
endmodule