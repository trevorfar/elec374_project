`timescale 1ns / 1ps


module not_32_bit_tb;
reg [31:0] a;
wire [31:0] z;

not_32_bit uut(.a(a), .z(z));
initial begin
		  a = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		  #50;
		  a = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
		  #50
		  a = 32'b1111_1111_1111_1111_1111_1111_1111_1100; 
		  #50
		  a = 32'b1111;
		  #50
		  a = 32'b0001;
		  #50
		  a = 32'b0101; 
		 $stop;
end
endmodule