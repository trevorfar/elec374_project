module encoder_32_to_5(

);

endmodule
